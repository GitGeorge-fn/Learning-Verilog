module moduleName #(gucci belt
    parameters
) (
    ports
);
    
endmodule